library ieee;
use ieee.std_logic_1164.all;

package char is
    function char_to_bits(signal char: character) return std_logic_vector;
    function bits_to_char(signal bits: std_logic_vector) return character;
end package;

package body char is

    function char_to_bits(signal char: in character)
    -- Converts a character to the ASCII binary representation
    return std_logic_vector is variable bits: std_logic_vector(7 downto 0);
    begin
        case char is
            when ' ' => bits := "00100000";
            when '!' => bits := "00100001";
            when '"' => bits := "00100010";
            when '#' => bits := "00100011";
            when '$' => bits := "00100100";
            -- when '%' => bits := "00100101";
            when '&' => bits := "00100110";
            when ''' => bits := "00100111";
            when '(' => bits := "00101000";
            when ')' => bits := "00101001";
            when '*' => bits := "00101010";
            when '+' => bits := "00101011";
            when ',' => bits := "00101100";
            when '-' => bits := "00101101";
            when '.' => bits := "00101110";
            when '/' => bits := "00101111";
            when '0' => bits := "00110000";
            when '1' => bits := "00110001";
            when '2' => bits := "00110010";
            when '3' => bits := "00110011";
            when '4' => bits := "00110100";
            when '5' => bits := "00110101";
            when '6' => bits := "00110110";
            when '7' => bits := "00110111";
            when '8' => bits := "00111000";
            when '9' => bits := "00111001";
            when ':' => bits := "00111010";
            when ';' => bits := "00111011";
            when '<' => bits := "00111100";
            when '=' => bits := "00111101";
            when '>' => bits := "00111110";
            when '?' => bits := "00111111";
            when '@' => bits := "01000000";
            when 'A' => bits := "01000001";
            when 'B' => bits := "01000010";
            when 'C' => bits := "01000011";
            when 'D' => bits := "01000100";
            when 'E' => bits := "01000101";
            when 'F' => bits := "01000110";
            when 'G' => bits := "01000111";
            when 'H' => bits := "01001000";
            when 'I' => bits := "01001001";
            when 'J' => bits := "01001010";
            when 'K' => bits := "01001011";
            when 'L' => bits := "01001100";
            when 'M' => bits := "01001101";
            when 'N' => bits := "01001110";
            when 'O' => bits := "01001111";
            when 'P' => bits := "01010000";
            when 'Q' => bits := "01010001";
            when 'R' => bits := "01010010";
            when 'S' => bits := "01010011";
            when 'T' => bits := "01010100";
            when 'U' => bits := "01010101";
            when 'V' => bits := "01010110";
            when 'W' => bits := "01010111";
            when 'X' => bits := "01011000";
            when 'Y' => bits := "01011001";
            when 'Z' => bits := "01011010";
            when '[' => bits := "01011011";
            when '\' => bits := "01011100";
            when ']' => bits := "01011101";
            when '^' => bits := "01011110";
            when '_' => bits := "01011111";
            when '`' => bits := "01100000";
            when 'a' => bits := "01100001";
            when 'b' => bits := "01100010";
            when 'c' => bits := "01100011";
            when 'd' => bits := "01100100";
            when 'e' => bits := "01100101";
            when 'f' => bits := "01100110";
            when 'g' => bits := "01100111";
            when 'h' => bits := "01101000";
            when 'i' => bits := "01101001";
            when 'j' => bits := "01101010";
            when 'k' => bits := "01101011";
            when 'l' => bits := "01101100";
            when 'm' => bits := "01101101";
            when 'n' => bits := "01101110";
            when 'o' => bits := "01101111";
            when 'p' => bits := "01110000";
            when 'q' => bits := "01110001";
            when 'r' => bits := "01110010";
            when 's' => bits := "01110011";
            when 't' => bits := "01110100";
            when 'u' => bits := "01110101";
            when 'v' => bits := "01110110";
            when 'w' => bits := "01110111";
            when 'x' => bits := "01111000";
            when 'y' => bits := "01111001";
            when 'z' => bits := "01111010";
            when '{' => bits := "01111011";
            when '|' => bits := "01111100";
            when '}' => bits := "01111101";
            when '~' => bits := "01111110";
            when others => bits := "11111111";
        end case;
        return bits;
    end char_to_bits;
    
    function bits_to_char(signal bits: in std_logic_vector(6 downto 0))
    -- Converts a custom BCD-like representation to the corresponding character
    return character is variable char: character;
    begin
        case bits is
            when "0000000" => char := ' '; when "1000000" => char := ' ';
            when "0000001" => char := 'a';
            when "0000010" => char := 'b';
            when "0000011" => char := 'c';
            when "0000100" => char := 'd';
            when "0000101" => char := 'e';
            when "0000110" => char := 'f';
            when "0000111" => char := 'g';
            when "0001000" => char := 'h';
            when "0001001" => char := 'i';
            when "0010000" => char := 'j';
            when "0010001" => char := 'k';
            when "0010010" => char := 'l';
            when "0010011" => char := 'm';
            when "0010100" => char := 'n';
            when "0010101" => char := 'o';
            when "0010110" => char := 'p';
            when "0010111" => char := 'q';
            when "0011000" => char := 'r';
            when "0011001" => char := 's';
            when "0100000" => char := 't';
            when "0100001" => char := 'u';
            when "0100010" => char := 'v';
            when "0100011" => char := 'w';
            when "0100100" => char := 'x';
            when "0100101" => char := 'y';
            when "0100110" => char := 'z';
            when "1000001" => char := 'A';
            when "1000010" => char := 'B';
            when "1000011" => char := 'C';
            when "1000100" => char := 'D';
            when "1000101" => char := 'E';
            when "1000110" => char := 'F';
            when "1000111" => char := 'G';
            when "1001000" => char := 'H';
            when "1001001" => char := 'I';
            when "1010000" => char := 'J';
            when "1010001" => char := 'K';
            when "1010010" => char := 'L';
            when "1010011" => char := 'M';
            when "1010100" => char := 'N';
            when "1010101" => char := 'O';
            when "1010110" => char := 'P';
            when "1010111" => char := 'Q';
            when "1011000" => char := 'R';
            when "1011001" => char := 'S';
            when "1100000" => char := 'T';
            when "1100001" => char := 'U';
            when "1100010" => char := 'V';
            when "1100011" => char := 'W';
            when "1100100" => char := 'X';
            when "1100101" => char := 'Y';
            when "1100110" => char := 'Z';
            when "0100111" => char := ','; when "1100111" => char := ',';
            when "0101000" => char := '.'; when "1101000" => char := '.';
            when "0101001" => char := '-'; when "1101001" => char := '-';
            when "0110000" => char := '0'; when "1110000" => char := '0';
            when "0110001" => char := '1'; when "1110001" => char := '1';
            when "0110010" => char := '2'; when "1110010" => char := '2';
            when "0110011" => char := '3'; when "1110011" => char := '3';
            when "0110100" => char := '4'; when "1110100" => char := '4';
            when "0110101" => char := '5'; when "1110101" => char := '5';
            when "0110110" => char := '6'; when "1110110" => char := '6';
            when "0110111" => char := '7'; when "1110111" => char := '7';
            when "0111000" => char := '8'; when "1111000" => char := '8';
            when "0111001" => char := '9'; when "1111001" => char := '9';
            when others => char := nul;
        end case;
        return char;
    end bits_to_char;

end char;
